module branch_control(
    input zero,
    input branch,
    output [31:0] result
);

